// module decoder with 5 inputes and 2n outputs
module decoder(
    input [4:0] a, en,
    output [31:0] y
    );
    always @(in) begin
        if (a) begin
            y = 32'b0
            case (a or en)
                5'b00000: y[0] = ;
                5'b00001: y[1] = ;
                5'b00010: y[2] = ;
                5'b00011: y[3] = ;
                5'b00100: y[4] = ;
                5'b00101: y[5] = ;
                5'b00110: y[6] = ;
                5'b00111: y[7] = ;
                5'b01000: y[8] = ;
                5'b01001: y[9] = ;
                5'b01010: y[10] = ;
                5'b01011: y[11] = ;
                5'b01100: y[12] = ;
                5'b01101: y[13] = ;
                5'b01110: y[14] = ;
                5'b01111: y[15] = ;
                5'b10000: y[16] = ;
                5'b10001: y[17] = ;
                5'b10010: y[18] = ;
                5'b10011: y[19] = ;
                5'b10100: y[20] = ;
                5'b10101: y[21] = ;
                5'b10110: y[22] = ;
                5'b10111: y[23] = ;
                5'b11000: y[24] = ;
                5'b11001: y[25] = ;
                5'b11010: y[26] = 0;
                5'b11011: y[27] = 0;
                5'b11100: y[28] = 0;
                5'b11101: y[29] = 0;
                5'b11110: y[30] = 0;
                5'b11111: y[31] = 0;
                default: 
            endcase
        end
    end
endmodule
